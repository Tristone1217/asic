this is a useful example
this is a useful example for linux command study
this is a useful example for my linux command study
useful example useful example  useful example useful example useful example useful example
