this is a example
this is a example for linux command study
this is a example for my linux command study
example example  example example example example
